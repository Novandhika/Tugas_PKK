`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/06/2022 04:20:37 PM
// Design Name: 
// Module Name: instr_mem
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module instr_mem(
	input			clk,
	input[31:0]		addr,
	output [31:0]	instr
	);
	
	reg[31:0]	out;
	assign instr = out;
	always@(posedge clk)
	begin
		case(addr)
			32'd0	:	out = 32'b000000000001_00000_000_00101_0010011;//ADDI rd = 5 , rs1 = 0, func3 = 0 , imm = 1
			32'd1	:	out = 32'b000000000101_00000_000_00110_0010011;//ADDI rd = 6 , rs1 = 0, func3 = 0 , imm = 5
			32'd2	:	out = 32'b111111111111_00000_000_00111_0010011;//ADDI rd = 7 , rs1 = 0, func3 = 0 , imm = -1
			32'd3	:	out = 32'b0_000000_00101_00101_000_0001_0_1100011;//BEQ imm = 2 , rs1 = 5 , rs2 = 5
			32'd4	:	out = 32'b000000000001_00000_000_11110_0010011;//ADDI rd = 30, func3 = 0 , imm = 1
			32'd5	:	out = 32'b0_000000_00000_00101_000_0000_0_1100011;//BEQ imm = 0 , rs1 = 5 , rs2 = 0
			32'd6	:	out = 32'b0_000000_00000_00101_001_0001_0_1100011;//BNE imm = 1 , rs1 = 5 , rs2 = 0
			32'd7	:	out = 32'b000000000001_00000_000_11110_0010011;//ADDI rd = 30, rs1 = 0, func3 = 0 , imm = 1
			32'd8	:	out = 32'b0_000000_00000_00000_001_0000_0_1100011;//BNE imm = 0, rs1 = 0, rs2 = 0
			32'd9	:	out = 32'b0_000000_00110_00111_100_0001_0_1100011;//BLT imm = 1, rs1 = 7, rs2 = 6
			32'd10	:	out = 32'b000000000001_00000_000_11110_0010011;//ADDI rd = 30, func3 = 0, rs1 = 0, imm = 1
			32'd11	:	out = 32'b0_000000_00111_00110_100_0000_0_1100011;//BLT imm = 0, rs1 = 6, rs2 = 7
			32'd12	:	out = 32'b0_000000_00111_00110_101_0001_0_1100011;//BGE imm = 1, rs1 = 6, rs2 = 7
			32'd13	:	out = 32'b000000000001_00000_000_11110_0010011;//ADDI rd = 30, rs1 = 0, funct3 = 0, imm = 1
			32'd14	:	out = 32'b0_000000_00000_00111_101_0000_0_1100011;//BGE imm = 0, rs1 = 7, rs2 = 0
			32'd15	:	out = 32'b0_000000_00111_00101_110_0001_0_1100011;//BLTU imm = 1, rs1 = 5, rs2 = 7
			32'd16	:	out = 32'b000000000001_00000_000_11111_0010011;//ADDI rd = 31, rs1 = 0, func3 = 0, imm = 1
			32'd17	:	out = 32'b000000000010_00000_000_11111_0010011;//ADDI rd = 31, rs1 = 0, func3 = 0, imm = 2
			32'd18	:	out = 32'b1_111111_00000_00000_110_1110_1_1100011;//BLTU imm = -4, rs1 = 0, rs2 = 0
			32'd19	:	out = 32'b0_000000_00110_00111_111_0001_0_1100011;//BGEU imm = 1 , rs1 = 7, rs2 = 6
			32'd20	:	out = 32'b000000000001_00000_000_11110_0010011;
			32'd21	:	out = 32'b000000000001_11110_000_11110_0010011;
			32'd22	:	out = 32'b0000000000000000000000000_0000000; 
			default: out = 32'd0; 
		endcase
	end
	

endmodule
